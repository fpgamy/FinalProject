module lazy_shit(what_i_want1, what_i_want2);
output [29:0] what_i_want1;
output [29:0] what_i_want2;
assign what_i_want1 = 50;
assign what_i_want2 = 350;
endmodule